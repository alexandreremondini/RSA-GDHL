library verilog;
use verilog.vl_types.all;
entity INV3_3B is
    port(
        A               : in     vl_logic;
        Q               : out    vl_logic
    );
end INV3_3B;
