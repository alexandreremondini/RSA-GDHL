library verilog;
use verilog.vl_types.all;
entity TIE0_3B is
    port(
        Q               : out    vl_logic
    );
end TIE0_3B;
