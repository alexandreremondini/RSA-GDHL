library verilog;
use verilog.vl_types.all;
entity ITP_V5 is
    port(
        PAD             : in     vl_logic;
        Y               : out    vl_logic
    );
end ITP_V5;
