library verilog;
use verilog.vl_types.all;
entity BUDD8P is
    port(
        A               : in     vl_logic;
        PAD             : out    vl_logic
    );
end BUDD8P;
