library verilog;
use verilog.vl_types.all;
entity U_FJK_P_SB_NO is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end U_FJK_P_SB_NO;
