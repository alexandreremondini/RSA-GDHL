library verilog;
use verilog.vl_types.all;
entity BU12SP_3B is
    port(
        A               : in     vl_logic;
        PAD             : out    vl_logic
    );
end BU12SP_3B;
