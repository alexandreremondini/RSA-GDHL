library verilog;
use verilog.vl_types.all;
entity AVDD5ALLP_3B is
    port(
        A               : in     vl_logic
    );
end AVDD5ALLP_3B;
