library verilog;
use verilog.vl_types.all;
entity DLY22 is
    port(
        A               : in     vl_logic;
        Q               : out    vl_logic
    );
end DLY22;
