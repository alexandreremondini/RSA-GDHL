library verilog;
use verilog.vl_types.all;
entity ARAILPROT5P is
end ARAILPROT5P;
