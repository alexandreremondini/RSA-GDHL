library verilog;
use verilog.vl_types.all;
entity DLY32 is
    port(
        A               : in     vl_logic;
        Q               : out    vl_logic
    );
end DLY32;
