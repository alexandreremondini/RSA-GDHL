library verilog;
use verilog.vl_types.all;
entity U_FD_P_RB_NO is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end U_FD_P_RB_NO;
