library verilog;
use verilog.vl_types.all;
entity DLY42 is
    port(
        A               : in     vl_logic;
        Q               : out    vl_logic
    );
end DLY42;
