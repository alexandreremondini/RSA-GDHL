library verilog;
use verilog.vl_types.all;
entity BU8SP_3B is
    port(
        A               : in     vl_logic;
        PAD             : out    vl_logic
    );
end BU8SP_3B;
