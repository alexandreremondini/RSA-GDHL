library verilog;
use verilog.vl_types.all;
entity VDD5ALLP_V5 is
    port(
        A               : inout  vl_logic
    );
end VDD5ALLP_V5;
