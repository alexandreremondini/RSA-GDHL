library verilog;
use verilog.vl_types.all;
entity BUDD4P_V5 is
    port(
        A               : in     vl_logic;
        PAD             : out    vl_logic
    );
end BUDD4P_V5;
