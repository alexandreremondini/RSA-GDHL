library verilog;
use verilog.vl_types.all;
entity DFF_UDP is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end DFF_UDP;
