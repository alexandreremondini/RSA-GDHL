library verilog;
use verilog.vl_types.all;
entity ICP_3B is
    port(
        PAD             : in     vl_logic;
        Y               : out    vl_logic
    );
end ICP_3B;
