library verilog;
use verilog.vl_types.all;
entity ITCK2P_V5 is
    port(
        PAD             : in     vl_logic;
        Y               : out    vl_logic
    );
end ITCK2P_V5;
