library verilog;
use verilog.vl_types.all;
entity CLKIN12_3B is
    port(
        A               : in     vl_logic;
        Q               : out    vl_logic
    );
end CLKIN12_3B;
