library verilog;
use verilog.vl_types.all;
entity ICCK4P_V5 is
    port(
        PAD             : in     vl_logic;
        Y               : out    vl_logic
    );
end ICCK4P_V5;
