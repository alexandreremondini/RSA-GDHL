library verilog;
use verilog.vl_types.all;
entity APRIOP_3B is
    port(
        PAD             : inout  vl_logic;
        Z               : inout  vl_logic
    );
end APRIOP_3B;
