library verilog;
use verilog.vl_types.all;
entity ICUP_V5 is
    port(
        PAD             : in     vl_logic;
        Y               : out    vl_logic
    );
end ICUP_V5;
