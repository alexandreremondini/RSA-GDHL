library verilog;
use verilog.vl_types.all;
entity GND3OP is
    port(
        A               : inout  vl_logic
    );
end GND3OP;
