library verilog;
use verilog.vl_types.all;
entity AGND5ALLP_3B is
    port(
        A               : in     vl_logic
    );
end AGND5ALLP_3B;
