library verilog;
use verilog.vl_types.all;
entity BUDU2P_V5 is
    port(
        A               : in     vl_logic;
        PAD             : out    vl_logic
    );
end BUDU2P_V5;
