library verilog;
use verilog.vl_types.all;
entity VDD3ALLP is
    port(
        A               : inout  vl_logic
    );
end VDD3ALLP;
