library verilog;
use verilog.vl_types.all;
entity GND5IP_V5 is
    port(
        A               : inout  vl_logic
    );
end GND5IP_V5;
