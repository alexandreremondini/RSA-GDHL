library verilog;
use verilog.vl_types.all;
entity DLY32_3B is
    port(
        A               : in     vl_logic;
        Q               : out    vl_logic
    );
end DLY32_3B;
