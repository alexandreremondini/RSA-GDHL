library verilog;
use verilog.vl_types.all;
entity ICDP_3B is
    port(
        PAD             : in     vl_logic;
        Y               : out    vl_logic
    );
end ICDP_3B;
