library verilog;
use verilog.vl_types.all;
entity TIE0 is
    port(
        Q               : out    vl_logic
    );
end TIE0;
