library verilog;
use verilog.vl_types.all;
entity LOGIC0_3B is
    port(
        Q               : out    vl_logic
    );
end LOGIC0_3B;
