library verilog;
use verilog.vl_types.all;
entity INV0 is
    port(
        A               : in     vl_logic;
        Q               : out    vl_logic
    );
end INV0;
