library verilog;
use verilog.vl_types.all;
entity BU16SMP_3B is
    port(
        A               : in     vl_logic;
        PAD             : out    vl_logic
    );
end BU16SMP_3B;
