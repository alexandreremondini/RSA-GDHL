library verilog;
use verilog.vl_types.all;
entity AVDD3ALLP is
    port(
        VDDA            : in     vl_logic
    );
end AVDD3ALLP;
