library verilog;
use verilog.vl_types.all;
entity ITCK8P_3B is
    port(
        PAD             : in     vl_logic;
        Y               : out    vl_logic
    );
end ITCK8P_3B;
