library verilog;
use verilog.vl_types.all;
entity U_MUX_3_2_INV is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end U_MUX_3_2_INV;
