library verilog;
use verilog.vl_types.all;
entity ICP_V5 is
    port(
        PAD             : in     vl_logic;
        Y               : out    vl_logic
    );
end ICP_V5;
