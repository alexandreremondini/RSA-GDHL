library verilog;
use verilog.vl_types.all;
entity ISDP_V5 is
    port(
        PAD             : in     vl_logic;
        Y               : out    vl_logic
    );
end ISDP_V5;
