library verilog;
use verilog.vl_types.all;
entity ISUP_V5 is
    port(
        PAD             : in     vl_logic;
        Y               : out    vl_logic
    );
end ISUP_V5;
