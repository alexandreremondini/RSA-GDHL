library verilog;
use verilog.vl_types.all;
entity GND3RP is
    port(
        A               : inout  vl_logic
    );
end GND3RP;
