library verilog;
use verilog.vl_types.all;
entity ARAILPROT3P is
end ARAILPROT3P;
