library verilog;
use verilog.vl_types.all;
entity LOGIC0 is
    port(
        Q               : out    vl_logic
    );
end LOGIC0;
