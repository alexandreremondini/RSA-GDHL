library verilog;
use verilog.vl_types.all;
entity ICCK4P is
    port(
        PAD             : in     vl_logic;
        Y               : out    vl_logic
    );
end ICCK4P;
