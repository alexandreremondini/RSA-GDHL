library verilog;
use verilog.vl_types.all;
entity TIELOW is
    port(
        Q               : out    vl_logic
    );
end TIELOW;
