library verilog;
use verilog.vl_types.all;
entity APRIOWP is
    port(
        Z               : inout  vl_logic;
        PAD             : inout  vl_logic
    );
end APRIOWP;
