library verilog;
use verilog.vl_types.all;
entity GND3RP_3B is
    port(
        A               : inout  vl_logic
    );
end GND3RP_3B;
