library verilog;
use verilog.vl_types.all;
entity BUF4_3B is
    port(
        A               : in     vl_logic;
        Q               : out    vl_logic
    );
end BUF4_3B;
