library verilog;
use verilog.vl_types.all;
entity BUDD4P_3B is
    port(
        A               : in     vl_logic;
        PAD             : out    vl_logic
    );
end BUDD4P_3B;
