library verilog;
use verilog.vl_types.all;
entity BU8SP is
    port(
        A               : in     vl_logic;
        PAD             : out    vl_logic
    );
end BU8SP;
