library verilog;
use verilog.vl_types.all;
entity BUFE10 is
    port(
        A               : in     vl_logic;
        E               : in     vl_logic;
        Q               : out    vl_logic
    );
end BUFE10;
