library verilog;
use verilog.vl_types.all;
entity TIEHIGH_3B is
    port(
        Q               : out    vl_logic
    );
end TIEHIGH_3B;
