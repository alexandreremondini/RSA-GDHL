library verilog;
use verilog.vl_types.all;
entity ICCK16P is
    port(
        PAD             : in     vl_logic;
        Y               : out    vl_logic
    );
end ICCK16P;
