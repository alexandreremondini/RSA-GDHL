library verilog;
use verilog.vl_types.all;
entity VDD3RP is
    port(
        A               : inout  vl_logic
    );
end VDD3RP;
