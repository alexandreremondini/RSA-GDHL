library verilog;
use verilog.vl_types.all;
entity RAILPROTP_3B is
end RAILPROTP_3B;
