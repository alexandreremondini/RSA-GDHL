library verilog;
use verilog.vl_types.all;
entity BUDU8P_3B is
    port(
        A               : in     vl_logic;
        PAD             : out    vl_logic
    );
end BUDU8P_3B;
