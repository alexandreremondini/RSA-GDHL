library verilog;
use verilog.vl_types.all;
entity TIE1_3B is
    port(
        Q               : out    vl_logic
    );
end TIE1_3B;
