library verilog;
use verilog.vl_types.all;
entity LOGIC1 is
    port(
        Q               : out    vl_logic
    );
end LOGIC1;
