library verilog;
use verilog.vl_types.all;
entity CLKIN1 is
    port(
        A               : in     vl_logic;
        Q               : out    vl_logic
    );
end CLKIN1;
