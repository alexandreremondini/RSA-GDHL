library verilog;
use verilog.vl_types.all;
entity TIEHIGH is
    port(
        Q               : out    vl_logic
    );
end TIEHIGH;
