library verilog;
use verilog.vl_types.all;
entity ISUP_3B is
    port(
        PAD             : in     vl_logic;
        Y               : out    vl_logic
    );
end ISUP_3B;
