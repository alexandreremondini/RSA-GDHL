library verilog;
use verilog.vl_types.all;
entity GND5OP_V5 is
    port(
        A               : inout  vl_logic
    );
end GND5OP_V5;
