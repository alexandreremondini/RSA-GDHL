library verilog;
use verilog.vl_types.all;
entity BUFE12 is
    port(
        A               : in     vl_logic;
        E               : in     vl_logic;
        Q               : out    vl_logic
    );
end BUFE12;
