library verilog;
use verilog.vl_types.all;
entity CLKBU15_3B is
    port(
        A               : in     vl_logic;
        Q               : out    vl_logic
    );
end CLKBU15_3B;
