library verilog;
use verilog.vl_types.all;
entity TIELOW_3B is
    port(
        Q               : out    vl_logic
    );
end TIELOW_3B;
