library verilog;
use verilog.vl_types.all;
entity VDD3OP is
    port(
        A               : inout  vl_logic
    );
end VDD3OP;
