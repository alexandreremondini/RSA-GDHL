library verilog;
use verilog.vl_types.all;
entity BUDU16P_3B is
    port(
        A               : in     vl_logic;
        PAD             : out    vl_logic
    );
end BUDU16P_3B;
