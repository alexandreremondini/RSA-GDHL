library verilog;
use verilog.vl_types.all;
entity BUSHD_3B is
    port(
        A               : inout  vl_logic
    );
end BUSHD_3B;
