library verilog;
use verilog.vl_types.all;
entity AVDD3ALLP_3B is
    port(
        A               : in     vl_logic
    );
end AVDD3ALLP_3B;
