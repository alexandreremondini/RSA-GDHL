library verilog;
use verilog.vl_types.all;
entity INV0_3B is
    port(
        A               : in     vl_logic;
        Q               : out    vl_logic
    );
end INV0_3B;
