library verilog;
use verilog.vl_types.all;
entity RAILPROTP is
end RAILPROTP;
