library verilog;
use verilog.vl_types.all;
entity BUDD24P is
    port(
        A               : in     vl_logic;
        PAD             : out    vl_logic
    );
end BUDD24P;
