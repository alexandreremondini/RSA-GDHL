library verilog;
use verilog.vl_types.all;
entity ARAILPROT3P_3B is
end ARAILPROT3P_3B;
