library verilog;
use verilog.vl_types.all;
entity U_dfsecp_Q is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end U_dfsecp_Q;
