library verilog;
use verilog.vl_types.all;
entity CBU1P_3B is
    port(
        A               : in     vl_logic;
        Y               : out    vl_logic
    );
end CBU1P_3B;
