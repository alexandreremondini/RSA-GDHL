library verilog;
use verilog.vl_types.all;
entity DLY12_3B is
    port(
        A               : in     vl_logic;
        Q               : out    vl_logic
    );
end DLY12_3B;
