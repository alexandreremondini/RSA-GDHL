library verilog;
use verilog.vl_types.all;
entity APRIO1K5P_3B is
    port(
        PAD             : inout  vl_logic;
        Z               : inout  vl_logic
    );
end APRIO1K5P_3B;
