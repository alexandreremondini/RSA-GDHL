library verilog;
use verilog.vl_types.all;
entity APRIOWP_3B is
    port(
        PAD             : inout  vl_logic;
        Z               : inout  vl_logic
    );
end APRIOWP_3B;
