library verilog;
use verilog.vl_types.all;
entity CBU1P_V5 is
    port(
        A               : in     vl_logic;
        Y               : out    vl_logic
    );
end CBU1P_V5;
