library verilog;
use verilog.vl_types.all;
entity VDD3OP_3B is
    port(
        A               : inout  vl_logic
    );
end VDD3OP_3B;
