library verilog;
use verilog.vl_types.all;
entity APRIO200P is
    port(
        Z               : inout  vl_logic;
        PAD             : inout  vl_logic
    );
end APRIO200P;
