library verilog;
use verilog.vl_types.all;
entity BUSHD is
    port(
        A               : inout  vl_logic
    );
end BUSHD;
