library verilog;
use verilog.vl_types.all;
entity RAILPROTP_V5 is
end RAILPROTP_V5;
