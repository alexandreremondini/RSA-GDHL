library verilog;
use verilog.vl_types.all;
entity BUF8_3B is
    port(
        A               : in     vl_logic;
        Q               : out    vl_logic
    );
end BUF8_3B;
