library verilog;
use verilog.vl_types.all;
entity ITDP_V5 is
    port(
        PAD             : in     vl_logic;
        Y               : out    vl_logic
    );
end ITDP_V5;
