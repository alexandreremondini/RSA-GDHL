library verilog;
use verilog.vl_types.all;
entity AVSUBP_3B is
    port(
        A               : in     vl_logic
    );
end AVSUBP_3B;
