library verilog;
use verilog.vl_types.all;
entity ISP_3B is
    port(
        PAD             : in     vl_logic;
        Y               : out    vl_logic
    );
end ISP_3B;
