library verilog;
use verilog.vl_types.all;
entity ISDP is
    port(
        PAD             : in     vl_logic;
        Y               : out    vl_logic
    );
end ISDP;
