library verilog;
use verilog.vl_types.all;
entity CLKIN0 is
    port(
        A               : in     vl_logic;
        Q               : out    vl_logic
    );
end CLKIN0;
