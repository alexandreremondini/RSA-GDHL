library verilog;
use verilog.vl_types.all;
entity APRIO1K5P is
    port(
        Z               : inout  vl_logic;
        PAD             : inout  vl_logic
    );
end APRIO1K5P;
