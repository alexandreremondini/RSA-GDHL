library verilog;
use verilog.vl_types.all;
entity BUF12_3B is
    port(
        A               : in     vl_logic;
        Q               : out    vl_logic
    );
end BUF12_3B;
