library verilog;
use verilog.vl_types.all;
entity ISP_V5 is
    port(
        PAD             : in     vl_logic;
        Y               : out    vl_logic
    );
end ISP_V5;
