library verilog;
use verilog.vl_types.all;
entity DLY42_3B is
    port(
        A               : in     vl_logic;
        Q               : out    vl_logic
    );
end DLY42_3B;
