library verilog;
use verilog.vl_types.all;
entity AGND5ALLP is
    port(
        VSSA            : in     vl_logic
    );
end AGND5ALLP;
