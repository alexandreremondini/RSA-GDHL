library verilog;
use verilog.vl_types.all;
entity AGND3ALLP_3B is
    port(
        A               : in     vl_logic
    );
end AGND3ALLP_3B;
