library verilog;
use verilog.vl_types.all;
entity VDD3IP_V5 is
    port(
        A               : inout  vl_logic
    );
end VDD3IP_V5;
