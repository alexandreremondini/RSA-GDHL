library verilog;
use verilog.vl_types.all;
entity GND3IP is
    port(
        A               : inout  vl_logic
    );
end GND3IP;
