library verilog;
use verilog.vl_types.all;
entity DLY22_3B is
    port(
        A               : in     vl_logic;
        Q               : out    vl_logic
    );
end DLY22_3B;
