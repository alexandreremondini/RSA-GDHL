library verilog;
use verilog.vl_types.all;
entity VSUBP_3B is
    port(
        A               : inout  vl_logic
    );
end VSUBP_3B;
