library verilog;
use verilog.vl_types.all;
entity TIE1 is
    port(
        Q               : out    vl_logic
    );
end TIE1;
