library verilog;
use verilog.vl_types.all;
entity MUX_UDP is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end MUX_UDP;
