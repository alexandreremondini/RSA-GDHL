library verilog;
use verilog.vl_types.all;
entity CBU1P is
    port(
        A               : in     vl_logic;
        Y               : out    vl_logic
    );
end CBU1P;
