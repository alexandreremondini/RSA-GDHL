library verilog;
use verilog.vl_types.all;
entity ICDP_V5 is
    port(
        PAD             : in     vl_logic;
        Y               : out    vl_logic
    );
end ICDP_V5;
