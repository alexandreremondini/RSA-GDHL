library verilog;
use verilog.vl_types.all;
entity BU12P_V5 is
    port(
        A               : in     vl_logic;
        PAD             : out    vl_logic
    );
end BU12P_V5;
