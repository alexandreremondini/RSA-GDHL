library verilog;
use verilog.vl_types.all;
entity APRIO50P_3B is
    port(
        PAD             : inout  vl_logic;
        Z               : inout  vl_logic
    );
end APRIO50P_3B;
