library verilog;
use verilog.vl_types.all;
entity AGND3ALLP is
    port(
        VSSA            : in     vl_logic
    );
end AGND3ALLP;
