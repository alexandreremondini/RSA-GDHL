library verilog;
use verilog.vl_types.all;
entity CLKBU12_3B is
    port(
        A               : in     vl_logic;
        Q               : out    vl_logic
    );
end CLKBU12_3B;
