library verilog;
use verilog.vl_types.all;
entity BUF12 is
    port(
        A               : in     vl_logic;
        Q               : out    vl_logic
    );
end BUF12;
