library verilog;
use verilog.vl_types.all;
entity ARAILPRO5P_3B is
end ARAILPRO5P_3B;
