library verilog;
use verilog.vl_types.all;
entity BUDD1P_V5 is
    port(
        A               : in     vl_logic;
        PAD             : out    vl_logic
    );
end BUDD1P_V5;
