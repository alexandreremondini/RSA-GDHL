library verilog;
use verilog.vl_types.all;
entity ITCK2P is
    port(
        PAD             : in     vl_logic;
        Y               : out    vl_logic
    );
end ITCK2P;
