library verilog;
use verilog.vl_types.all;
entity LATCH_UDP is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end LATCH_UDP;
