library verilog;
use verilog.vl_types.all;
entity BU4SMP is
    port(
        A               : in     vl_logic;
        PAD             : out    vl_logic
    );
end BU4SMP;
