library verilog;
use verilog.vl_types.all;
entity AVDD5ALLP is
    port(
        VDDA            : in     vl_logic
    );
end AVDD5ALLP;
