library verilog;
use verilog.vl_types.all;
entity BU24SP_3B is
    port(
        A               : in     vl_logic;
        PAD             : out    vl_logic
    );
end BU24SP_3B;
