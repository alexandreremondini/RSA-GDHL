library verilog;
use verilog.vl_types.all;
entity ITCK16P_3B is
    port(
        PAD             : in     vl_logic;
        Y               : out    vl_logic
    );
end ITCK16P_3B;
