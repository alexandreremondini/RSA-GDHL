library verilog;
use verilog.vl_types.all;
entity LOGIC1_3B is
    port(
        Q               : out    vl_logic
    );
end LOGIC1_3B;
