library verilog;
use verilog.vl_types.all;
entity CLKBU6_3B is
    port(
        A               : in     vl_logic;
        Q               : out    vl_logic
    );
end CLKBU6_3B;
